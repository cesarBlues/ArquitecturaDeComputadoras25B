// https://github.com/cesarBlues
module _and
(
	input wire entradaA,
	input wire entradaB,
	output wire salidaC
);

	assign salidaC = entradaA & entradaB;

endmodule
